module adma_tx_sched
#(
    
) (
    
);
    
endmodule
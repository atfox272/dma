module adma_chn_arb
#(
    
) (
    
);
    
endmodule
module adma_wr_host
#(
    
) (
    
);
    
endmodule
module adma_chn_man
#(
    
) (
    
);
    
endmodule
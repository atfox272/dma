module adma_rd_host
#(
    
) (
    
);
    
endmodule
module adma_chn_buf
#(
    
) (
    
);
    
endmodule
module adma_data_buf
#(
    
) (
    
);
    
endmodule